mg45@ecegrid-thin2.ecn.purdue.edu.8848:1521110835